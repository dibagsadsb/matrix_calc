// ����ģ�飺�������ϵͳ
// ���ܣ����Ͽ��� FSM���������ʾ��LED ״ָ̬ʾ���Լ� UART �ӿ�
module matrix_calc_top(
    input clk,               // ϵͳʱ��
    input rst_n,             // ��λ�źţ�����Ч
    input [3:0] dip_switch,  // DIP ���أ�����ģʽѡ��
    input button_confirm,    // ����ȷ������
    input uart_rx,           // UART ���ն˿�
    output uart_tx,          // UART ���Ͷ˿�
    output [7:0] leds,       // LED ״ָ̬ʾ
    output [6:0] seg_display // 7 ���������ʾ
);
 
    // �ڲ��ź�
    wire [3:0] state;        // ��ǰ״̬��״̬����Ϊ4λ��
    wire start_calc;         // FSM �����Ŀ�ʼ�����ź�
    wire calc_done;          // ������ɱ�־
    wire error_flag;         // ϵͳ�����־
    wire [3:0] op_type;      // ���������ź�
    wire countdown_done;     // ����ʱ����ź�
    wire start_countdown;    // ��������ʱ�ź�

    // ���� FSM ģ��
    controller_fsm u_ctrl (
        .clk(clk), 
        .rst_n(rst_n),
        .button(button_confirm),  // ��������
        .mode_sel(dip_switch),    // ģʽѡ��
        .calc_done(calc_done),    // �����������
        .error_in(error_flag),    // ��������
        .countdown_done(countdown_done),  // ����ʱ�������
        .state(state),            // �����ǰ״̬
        .start_calc(start_calc),  // �����ʼ�����ź�
        .op_type(op_type),        // �����������
        .error_led(leds[7]),     // ����LED��������
        .start_countdown(start_countdown) // �����������ʱ
    );

    // �������ʾģ��
    seg_display u_seg (
        .clk(clk),
        .state(state),           // ����״̬��ʾ��Ӧ��Ϣ
        .op_type(op_type),       // ������������
        .seg(seg_display)
    );

    // LED ָʾģ��
    led_status u_led (
        .state(state),           // ����״̬������Ӧ LED
        .leds(leds[6:0])         // ֻ����ǰ7��LED��LED7��FSM��������
    );

    // ����ģ�飨UART���洢�����㣩B �� C ʵ��
    // ������Ҫ���� calc_done, error_flag, countdown_done ���ź�

endmodule