// LED ״̬��ʾģ�飨�����棩
// ���ܣ����� FSM ״̬������Ӧ LED ָʾϵͳ״̬
module led_status(
    input [3:0] state,    // FSM ״̬���루4λ��
    output reg [7:0] leds // LED �����ÿλ��Ӧһ��״̬
);

    always @(*) begin
        leds = 8'b0; // Ĭ������ LED Ϩ��
        case(state)
            4'd0: leds[0] = 1'b1; // S0_IDLE ����״̬������ LED0
            4'd1: leds[1] = 1'b1; // S1_MENU �˵�״̬������ LED1
            4'd2: leds[2] = 1'b1; // S2_INPUT �û����룬���� LED2
            4'd3: leds[3] = 1'b1; // S3_GEN ���ɾ��󣬵��� LED3
            4'd4: leds[4] = 1'b1; // S4_DISPLAY ��ʾ��������� LED4
            4'd5: leds[5] = 1'b1; // S5_COMPUTE ����ִ�У����� LED5
            4'd6: leds[7] = 1'b1; // S6_ERROR ϵͳ���󣬵��� LED7
            4'd7: leds[6] = 1'b1; // S7_STORE �洢���󣬵��� LED6
            4'd8: leds[3] = 1'b1; // S8_SELECT ѡ�������������LED3��������أ�
            4'd9: leds[2] = 1'b1; // S9_WAIT ����ʱ�ȴ�������LED2��������أ�
            default: leds = 8'b0;  // δ����״̬ȫ��
        endcase
    end

endmodule