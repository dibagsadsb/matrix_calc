// ����ģ�飺��״̬�� FSM�������󵹼�ʱ��
module controller_fsm(
    input clk,              // ϵͳʱ��
    input rst_n,            // �첽��λ������Ч
    input button,           // ����ȷ��
    input [3:0] mode_sel,   // ģʽѡ��
    input calc_done,        // ��������ź�
    input error_in,         // ��������
    input countdown_done,   // ����������ʱ����ź�
    output reg [3:0] state, // ��ǰ״̬
    output reg start_calc,  // ���������ź�
    output reg [3:0] op_type, // ��ǰ��������
    output reg error_led,   // ����ָʾ LED
    output reg start_countdown // ��������������ʱ�ź�
);

    // ״̬���루���ֲ��䣩
    parameter S0_IDLE       = 4'd0,
              S1_MENU       = 4'd1,
              S2_INPUT      = 4'd2,
              S3_GEN        = 4'd3,
              S4_DISPLAY    = 4'd4,
              S5_COMPUTE    = 4'd5,
              S6_ERROR      = 4'd6,
              S7_STORE      = 4'd7,
              S8_SELECT     = 4'd8,
              S9_WAIT       = 4'd9;

    reg [3:0] next_state;

    // ״̬�Ĵ������£����ֲ��䣩
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            state <= S0_IDLE;
        else
            state <= next_state;
    end

    // ----------------------------
    // ��һ״̬�߼����ؼ��޸ģ�
    // ----------------------------
    always @(*) begin
        next_state = state;
        case(state)
            S0_IDLE: next_state = S1_MENU;
            S1_MENU: begin
                if(button) begin
                    case(mode_sel)
                        4'b0001: next_state = S2_INPUT;
                        4'b0010: next_state = S3_GEN;
                        4'b0100: next_state = S4_DISPLAY;
                        4'b1000: next_state = S8_SELECT; // �����Ƚ���ѡ�������
                        default: next_state = S1_MENU;
                    endcase
                end
            end
            
            S2_INPUT:  next_state = S7_STORE;
            S7_STORE:  next_state = S1_MENU; // �洢��ɻز˵�
            
            S8_SELECT: begin
                if (error_in) 
                    next_state = S9_WAIT;    // ѡ�������뵹��ʱ
                else 
                    next_state = S5_COMPUTE; // ѡ����ȷ��ʼ����
            end
            
            S3_GEN:    next_state = S1_MENU;
            S4_DISPLAY: next_state = S1_MENU;
            
            S5_COMPUTE: begin
                if (error_in)
                    next_state = S9_WAIT;    // ���������뵹��ʱ
                else if (calc_done)
                    next_state = S4_DISPLAY; // ���������ʾ���
                else
                    next_state = S5_COMPUTE;
            end
            
            S6_ERROR:  next_state = S9_WAIT; // ����״ֱ̬�ӽ��뵹��ʱ
            
            S9_WAIT: begin
                if (button) 
                    next_state = S8_SELECT;  // ����ʱ�ڰ���������ѡ�������
                else if (countdown_done)
                    next_state = S1_MENU;    // ����ʱ�������ز˵�
                else
                    next_state = S9_WAIT;    // ��������ʱ
            end
            
            default:   next_state = S1_MENU;
        endcase
    end

    // ----------------------------
    // ����߼����޸ģ�
    // ----------------------------
    always @(*) begin
        start_calc = (state == S5_COMPUTE);
        error_led  = (state == S6_ERROR) || (state == S9_WAIT); // ����͵���ʱ����LED
        start_countdown = (state == S9_WAIT); // ��������ʱ
        
        // �����������
        if (state == S8_SELECT || state == S9_WAIT)
            op_type = {1'b0, mode_sel[2:0]}; // ѡ��͵���ʱ�ڼ䱣�ֲ�������
        else
            op_type = 4'd0;
    end

endmodule