// �߶��������ʾģ�飨֧������������ʾ��
module seg_display(
    input clk,               // ϵͳʱ��
    input [3:0] state,       // FSM ״̬����
    input [3:0] op_type,     // ������������������
    output reg [6:0] seg     // �߶�����������a-g��
);

    // ----------------------------
    // ����ʱ�����Ĵ���
    // ----------------------------
    reg [25:0] clk_count;    // ʱ�Ӽ��������ڲ��� 1 ����ģ����� 100 MHz��
    reg [3:0] sec_count;     // �������֧�� 0~9 �뵹��ʱ��

    always @(posedge clk) begin
        if(state == 4'd9) begin
            if(clk_count >= 100_000_000 - 1) begin
                clk_count <= 0;
                if(sec_count != 0)
                    sec_count <= sec_count - 1;
            end else begin
                clk_count <= clk_count + 1;
            end
        end else begin
            clk_count <= 0;
            sec_count <= 4'd9;
        end
    end

    // ----------------------------
    // �������ʾ�߼����ؼ��޸ģ�
    // ----------------------------
    always @(*) begin
        if(state == 4'd9) begin
            // �ȴ�״̬��ʾ����ʱ����
            case(sec_count)
                4'd9: seg = 7'b0001110; // 9
                4'd8: seg = 7'b0000000; // 8
                4'd7: seg = 7'b0000110; // 7
                4'd6: seg = 7'b0100000; // 6
                4'd5: seg = 7'b0010010; // 5
                4'd4: seg = 7'b0110000; // 4
                4'd3: seg = 7'b0000110; // 3
                4'd2: seg = 7'b0010010; // 2
                4'd1: seg = 7'b1001111; // 1
                4'd0: seg = 7'b0000001; // 0
                default: seg = 7'b1111111;
            endcase
        end else if(state == 4'd8) begin
            // ��������ѡ�������״̬��ʾ��������
            case(op_type)
                4'b0001: seg = 7'b0000111; // T - ת��
                4'b0010: seg = 7'b0001000; // A - �ӷ�  
                4'b0100: seg = 7'b0000011; // B - �����˷�
                4'b1000: seg = 7'b1000110; // C - ����˷�
                default: seg = 7'b1111111; // Ĭ��ȫ��
            endcase
        end else begin
            // ����״̬����FSM״̬��ʾ�ַ�
            case(state)
                4'd0: seg = 7'b1111110; // I - ���У�S0_IDLE��
                4'd1: seg = 7'b0110000; // n - �˵���S1_MENU��
                4'd2: seg = 7'b1000000; // A - �û����루S2_INPUT��
                4'd3: seg = 7'b0001000; // G - ���ɾ���S3_GEN��
                4'd4: seg = 7'b0001001; // d - ��ʾ�����S4_DISPLAY��
                4'd5: seg = 7'b0000010; // C - ����ִ�У�S5_COMPUTE��
                4'd6: seg = 7'b0000110; // E - ϵͳ����S6_ERROR��
                4'd7: seg = 7'b0100001; // S7_STORE - �洢
                default: seg = 7'b1111111; // ����״̬ȫ��
            endcase
        end
    end

endmodule