// File: defs.vh
// ������㹤�̵�ȫ�ֲ�������
// ������ʹ�ñ��ļ������� .v �ļ��м��룺`include "defs.vh"

// �������ߴ磨��/�У�
`define MATRIX_MAX_SIZE           4       // ֧�� 4x4 ����
`define MATRIX_WIDTH              8       // �����ÿ��Ԫ���� 8-bit ����

// UART ����
`define UART_BAUD                 115200  // ���ڲ�����
`define CLK_FREQ                  100_000_000  // FPGA ������ʱ�� 100MHz

// ========== ״̬������ ==========���ؼ��޸ģ�
`define STATE_WIDTH               4       // ������״̬λ����
`define STATE_IDLE                4'd0    // ����
`define STATE_MENU                4'd1    // �˵���ʾ
`define STATE_INPUT               4'd2    // �û�����
`define STATE_GENERATE            4'd3    // �������Ծ���
`define STATE_DISPLAY             4'd4    // ��ʾ���
`define STATE_COMPUTE             4'd5    // ����ִ��
`define STATE_ERROR               4'd6    // ϵͳ����
`define STATE_STORE               4'd7    // �洢����
`define STATE_SELECT              4'd8    // ѡ�������
`define STATE_WAIT                4'd9    // ����ʱ�ȴ�

// ��ز������壨����չ��
`define DEBOUNCE_DELAY            20_000_000   // ����ȥ���ӳ�

// UART ��ز���
`define UART_START_BIT            1'b0
`define UART_STOP_BIT             1'b1
`define UART_DATA_BITS            8
`define UART_PARITY_ENABLE        0